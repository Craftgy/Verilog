module ptosda(rst,sclk,ack,scl,sda,data);

endmodule