module seqdet (
    ports
);
    
endmodule