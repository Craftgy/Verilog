`timescale 1ns/1ns
`define halfperiod 20

module t;
reg clk,rst;
reg[]
endmodule