`timescale 1ns/1ns
`define timeslice 100
module EEPROM(scl,sda);

endmodule