`timescale 1ns/1ns
module EEPROM();

endmodule