module seqdet (
    x,z,clk,rst
);
input x,clk,rst;
output z;
reg [2:0] state;

endmodule