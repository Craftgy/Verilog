`include "/Users/craft/资料/verilog_study/test.php/时序逻辑/状态机/fsm.v"
`timescale 1ns/1ns
module test