module seqdet (
    x,z,clk,rst
);
input 
endmodule