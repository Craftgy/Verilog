module out16hi(scl,sda,outh);

endmodule