module ptosda(rst,sclk,ack,scl,sda,data);
input sclk,rst;
inpu

endmodule