module seqdet (
    x,z,
);
    
endmodule