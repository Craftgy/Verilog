module pto();

endmodule