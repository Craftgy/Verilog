module out16hi();

endmodule