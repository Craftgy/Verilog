module ptosda();

endmodule