module seqdet (
    x,z,clk,rst
);
input x,clk
endmodule