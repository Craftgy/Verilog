module ptosda(rst,sclk,ack,scl,sda,);

endmodule