`timescale 1ns/1ns
`define halfperiod 50
module sigdata(rst,sclk,data,ask_for);

endmodule
