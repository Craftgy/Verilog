module out16hi(scl,sda,out);

endmodule