`timescale 1ns/1ns
module EEPROM_WR(SDA,SCL,ACK,RESET,CLK);

endmodule