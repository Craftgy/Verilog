module seqdet (
    
);
    
endmodule