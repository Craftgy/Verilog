module ptosda(rst,clk);

endmodule