`timescale 1ns/1ns
`define halfperiod 50
module si();

endmodule
