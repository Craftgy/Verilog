module ptosda(rst,sclk,ack,scl,sda,data);
input sclk,rst;
input [3:0]

endmodule