module out16hi(scl,sda,outhigh);
input scl,sda
endmodule