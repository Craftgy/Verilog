module out();

endmodule