module Se (
    ports
);
    
endmodule