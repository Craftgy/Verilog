module out16hi(scl,sda,outhigh);
input scl,sda;
output [15:0] outhigh;

endmodule