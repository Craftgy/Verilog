module out16hi(scl,sda,outhigh);

endmodule