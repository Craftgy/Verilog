module seqdet (
    x,z,clk,rst
);
    
endmodule