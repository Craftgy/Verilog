module ptosda(rst,sclk,);

endmodule