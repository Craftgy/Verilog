module seqdet (
    x,z,clk,rst
);
input x,clk,rst;
output z;

endmodule